netcdf file_util_test_data {
dimensions:
	x = 4 ;
	y = 3 ;
	z = 1 ;
variables:
	double var1(x) ;
	double var2(y) ;
	double table(y, x, z) ;
data:

 var1 = 1.0, 2.0, 3.0, 4.0 ;

 var2 = 10.0, 20.0, 30.0 ;

 table =
  1.0,
  2.0,
  3.0,
  4.0,
  10.0,
  20.0,
  30.0,
  40.0,
  100.0,
  200.0,
  300.0,
  400.0 ;
}
